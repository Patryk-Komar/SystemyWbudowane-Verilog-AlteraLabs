module binary_search (
	);
endmodule