module word_with_space (
	output [0:6] HEX0,HEX1,HEX2,HEX3,HEX4,HEX5);
	assign HEX0 = 7'b0100100;
	assign HEX1 = 7'b0110000;
	assign HEX2 = 7'b1001111;
	assign HEX3 = 7'b0011000;
	assign HEX4 = 7'b1111111;
	assign HEX5 = 7'b1111111;
endmodule