module liczba_bitow (
	input ,
	output);
	
endmodule